
module loader0 (
	noe_in);	

	input		noe_in;
endmodule
