module serial_loader();



	loader0 u0 (
		.noe_in (0)  // noe_in.noe
	);



endmodule 